`ifndef APB_MASTER_DEF

`define APB_MASTER_DEF

`define INACTIVE    2'b00
`define SETUP   	2'b01
`define ACTIVE  	2'b10

`define WRITE   	1'b1
`define READ    	1'b0

`endif

