`ifndef UART_DEF

`define UART_DEF

`define IDLE          3'b000
`define START         3'b001
`define DATA_BITS     3'b010
`define STOP          3'b011
`define CLEANUP       3'b100

`endif